            10'd0: sample = -10;
            10'd1, 10'd2: sample = -9;
            10'd3, 10'd4, 10'd5, 10'd6, 10'd7: sample = -8;
            10'd8, 10'd9, 10'd10, 10'd11, 10'd12, 10'd13, 10'd14, 10'd15, 10'd16, 10'd17, 10'd18: sample = -7;
            10'd19, 10'd20, 10'd21, 10'd22, 10'd23, 10'd24, 10'd25, 10'd26, 10'd27, 10'd28, 10'd29, 10'd30, 10'd31, 10'd32, 10'd33, 10'd34, 10'd35, 10'd36, 10'd37, 10'd38, 10'd39: sample = -6;
            10'd40, 10'd41, 10'd42, 10'd43, 10'd44, 10'd45, 10'd46, 10'd47, 10'd48, 10'd49, 10'd50, 10'd51, 10'd52, 10'd53, 10'd54, 10'd55, 10'd56, 10'd57, 10'd58, 10'd59, 10'd60, 10'd61, 10'd62, 10'd63, 10'd64, 10'd65, 10'd66, 10'd67, 10'd68, 10'd69, 10'd70, 10'd71, 10'd72, 10'd73, 10'd74, 10'd75, 10'd76: sample = -5;
            10'd77, 10'd78, 10'd79, 10'd80, 10'd81, 10'd82, 10'd83, 10'd84, 10'd85, 10'd86, 10'd87, 10'd88, 10'd89, 10'd90, 10'd91, 10'd92, 10'd93, 10'd94, 10'd95, 10'd96, 10'd97, 10'd98, 10'd99, 10'd100, 10'd101, 10'd102, 10'd103, 10'd104, 10'd105, 10'd106, 10'd107, 10'd108, 10'd109, 10'd110, 10'd111, 10'd112, 10'd113, 10'd114, 10'd115, 10'd116, 10'd117, 10'd118, 10'd119, 10'd120, 10'd121, 10'd122, 10'd123, 10'd124, 10'd125, 10'd126, 10'd127, 10'd128, 10'd129, 10'd130, 10'd131, 10'd132, 10'd133: sample = -4;
            10'd134, 10'd135, 10'd136, 10'd137, 10'd138, 10'd139, 10'd140, 10'd141, 10'd142, 10'd143, 10'd144, 10'd145, 10'd146, 10'd147, 10'd148, 10'd149, 10'd150, 10'd151, 10'd152, 10'd153, 10'd154, 10'd155, 10'd156, 10'd157, 10'd158, 10'd159, 10'd160, 10'd161, 10'd162, 10'd163, 10'd164, 10'd165, 10'd166, 10'd167, 10'd168, 10'd169, 10'd170, 10'd171, 10'd172, 10'd173, 10'd174, 10'd175, 10'd176, 10'd177, 10'd178, 10'd179, 10'd180, 10'd181, 10'd182, 10'd183, 10'd184, 10'd185, 10'd186, 10'd187, 10'd188, 10'd189, 10'd190, 10'd191, 10'd192, 10'd193, 10'd194, 10'd195, 10'd196, 10'd197, 10'd198, 10'd199, 10'd200, 10'd201, 10'd202, 10'd203, 10'd204, 10'd205, 10'd206, 10'd207, 10'd208, 10'd209, 10'd210, 10'd211, 10'd212, 10'd213: sample = -3;
            10'd214, 10'd215, 10'd216, 10'd217, 10'd218, 10'd219, 10'd220, 10'd221, 10'd222, 10'd223, 10'd224, 10'd225, 10'd226, 10'd227, 10'd228, 10'd229, 10'd230, 10'd231, 10'd232, 10'd233, 10'd234, 10'd235, 10'd236, 10'd237, 10'd238, 10'd239, 10'd240, 10'd241, 10'd242, 10'd243, 10'd244, 10'd245, 10'd246, 10'd247, 10'd248, 10'd249, 10'd250, 10'd251, 10'd252, 10'd253, 10'd254, 10'd255, 10'd256, 10'd257, 10'd258, 10'd259, 10'd260, 10'd261, 10'd262, 10'd263, 10'd264, 10'd265, 10'd266, 10'd267, 10'd268, 10'd269, 10'd270, 10'd271, 10'd272, 10'd273, 10'd274, 10'd275, 10'd276, 10'd277, 10'd278, 10'd279, 10'd280, 10'd281, 10'd282, 10'd283, 10'd284, 10'd285, 10'd286, 10'd287, 10'd288, 10'd289, 10'd290, 10'd291, 10'd292, 10'd293, 10'd294, 10'd295, 10'd296, 10'd297, 10'd298, 10'd299, 10'd300, 10'd301, 10'd302, 10'd303, 10'd304, 10'd305, 10'd306, 10'd307, 10'd308, 10'd309, 10'd310, 10'd311, 10'd312, 10'd313, 10'd314, 10'd315, 10'd316: sample = -2;
            10'd317, 10'd318, 10'd319, 10'd320, 10'd321, 10'd322, 10'd323, 10'd324, 10'd325, 10'd326, 10'd327, 10'd328, 10'd329, 10'd330, 10'd331, 10'd332, 10'd333, 10'd334, 10'd335, 10'd336, 10'd337, 10'd338, 10'd339, 10'd340, 10'd341, 10'd342, 10'd343, 10'd344, 10'd345, 10'd346, 10'd347, 10'd348, 10'd349, 10'd350, 10'd351, 10'd352, 10'd353, 10'd354, 10'd355, 10'd356, 10'd357, 10'd358, 10'd359, 10'd360, 10'd361, 10'd362, 10'd363, 10'd364, 10'd365, 10'd366, 10'd367, 10'd368, 10'd369, 10'd370, 10'd371, 10'd372, 10'd373, 10'd374, 10'd375, 10'd376, 10'd377, 10'd378, 10'd379, 10'd380, 10'd381, 10'd382, 10'd383, 10'd384, 10'd385, 10'd386, 10'd387, 10'd388, 10'd389, 10'd390, 10'd391, 10'd392, 10'd393, 10'd394, 10'd395, 10'd396, 10'd397, 10'd398, 10'd399, 10'd400, 10'd401, 10'd402, 10'd403, 10'd404, 10'd405, 10'd406, 10'd407, 10'd408, 10'd409, 10'd410, 10'd411, 10'd412, 10'd413, 10'd414, 10'd415, 10'd416, 10'd417, 10'd418, 10'd419, 10'd420, 10'd421, 10'd422, 10'd423, 10'd424, 10'd425, 10'd426, 10'd427, 10'd428, 10'd429, 10'd430, 10'd431, 10'd432, 10'd433, 10'd434, 10'd435: sample = -1;
            10'd436, 10'd437, 10'd438, 10'd439, 10'd440, 10'd441, 10'd442, 10'd443, 10'd444, 10'd445, 10'd446, 10'd447, 10'd448, 10'd449, 10'd450, 10'd451, 10'd452, 10'd453, 10'd454, 10'd455, 10'd456, 10'd457, 10'd458, 10'd459, 10'd460, 10'd461, 10'd462, 10'd463, 10'd464, 10'd465, 10'd466, 10'd467, 10'd468, 10'd469, 10'd470, 10'd471, 10'd472, 10'd473, 10'd474, 10'd475, 10'd476, 10'd477, 10'd478, 10'd479, 10'd480, 10'd481, 10'd482, 10'd483, 10'd484, 10'd485, 10'd486, 10'd487, 10'd488, 10'd489, 10'd490, 10'd491, 10'd492, 10'd493, 10'd494, 10'd495, 10'd496, 10'd497, 10'd498, 10'd499, 10'd500, 10'd501, 10'd502, 10'd503, 10'd504, 10'd505, 10'd506, 10'd507, 10'd508, 10'd509, 10'd510, 10'd511, 10'd512, 10'd513, 10'd514, 10'd515, 10'd516, 10'd517, 10'd518, 10'd519, 10'd520, 10'd521, 10'd522, 10'd523, 10'd524, 10'd525, 10'd526, 10'd527, 10'd528, 10'd529, 10'd530, 10'd531, 10'd532, 10'd533, 10'd534, 10'd535, 10'd536, 10'd537, 10'd538, 10'd539, 10'd540, 10'd541, 10'd542, 10'd543, 10'd544, 10'd545, 10'd546, 10'd547, 10'd548, 10'd549, 10'd550, 10'd551, 10'd552, 10'd553, 10'd554, 10'd555, 10'd556, 10'd557, 10'd558, 10'd559, 10'd560: sample = 0;
            10'd561, 10'd562, 10'd563, 10'd564, 10'd565, 10'd566, 10'd567, 10'd568, 10'd569, 10'd570, 10'd571, 10'd572, 10'd573, 10'd574, 10'd575, 10'd576, 10'd577, 10'd578, 10'd579, 10'd580, 10'd581, 10'd582, 10'd583, 10'd584, 10'd585, 10'd586, 10'd587, 10'd588, 10'd589, 10'd590, 10'd591, 10'd592, 10'd593, 10'd594, 10'd595, 10'd596, 10'd597, 10'd598, 10'd599, 10'd600, 10'd601, 10'd602, 10'd603, 10'd604, 10'd605, 10'd606, 10'd607, 10'd608, 10'd609, 10'd610, 10'd611, 10'd612, 10'd613, 10'd614, 10'd615, 10'd616, 10'd617, 10'd618, 10'd619, 10'd620, 10'd621, 10'd622, 10'd623, 10'd624, 10'd625, 10'd626, 10'd627, 10'd628, 10'd629, 10'd630, 10'd631, 10'd632, 10'd633, 10'd634, 10'd635, 10'd636, 10'd637, 10'd638, 10'd639, 10'd640, 10'd641, 10'd642, 10'd643, 10'd644, 10'd645, 10'd646, 10'd647, 10'd648, 10'd649, 10'd650, 10'd651, 10'd652, 10'd653, 10'd654, 10'd655, 10'd656, 10'd657, 10'd658, 10'd659, 10'd660, 10'd661, 10'd662, 10'd663, 10'd664, 10'd665, 10'd666, 10'd667, 10'd668, 10'd669, 10'd670, 10'd671, 10'd672, 10'd673, 10'd674, 10'd675, 10'd676, 10'd677, 10'd678, 10'd679: sample = 1;
            10'd680, 10'd681, 10'd682, 10'd683, 10'd684, 10'd685, 10'd686, 10'd687, 10'd688, 10'd689, 10'd690, 10'd691, 10'd692, 10'd693, 10'd694, 10'd695, 10'd696, 10'd697, 10'd698, 10'd699, 10'd700, 10'd701, 10'd702, 10'd703, 10'd704, 10'd705, 10'd706, 10'd707, 10'd708, 10'd709, 10'd710, 10'd711, 10'd712, 10'd713, 10'd714, 10'd715, 10'd716, 10'd717, 10'd718, 10'd719, 10'd720, 10'd721, 10'd722, 10'd723, 10'd724, 10'd725, 10'd726, 10'd727, 10'd728, 10'd729, 10'd730, 10'd731, 10'd732, 10'd733, 10'd734, 10'd735, 10'd736, 10'd737, 10'd738, 10'd739, 10'd740, 10'd741, 10'd742, 10'd743, 10'd744, 10'd745, 10'd746, 10'd747, 10'd748, 10'd749, 10'd750, 10'd751, 10'd752, 10'd753, 10'd754, 10'd755, 10'd756, 10'd757, 10'd758, 10'd759, 10'd760, 10'd761, 10'd762, 10'd763, 10'd764, 10'd765, 10'd766, 10'd767, 10'd768, 10'd769, 10'd770, 10'd771, 10'd772, 10'd773, 10'd774, 10'd775, 10'd776, 10'd777, 10'd778, 10'd779, 10'd780, 10'd781, 10'd782: sample = 2;
            10'd783, 10'd784, 10'd785, 10'd786, 10'd787, 10'd788, 10'd789, 10'd790, 10'd791, 10'd792, 10'd793, 10'd794, 10'd795, 10'd796, 10'd797, 10'd798, 10'd799, 10'd800, 10'd801, 10'd802, 10'd803, 10'd804, 10'd805, 10'd806, 10'd807, 10'd808, 10'd809, 10'd810, 10'd811, 10'd812, 10'd813, 10'd814, 10'd815, 10'd816, 10'd817, 10'd818, 10'd819, 10'd820, 10'd821, 10'd822, 10'd823, 10'd824, 10'd825, 10'd826, 10'd827, 10'd828, 10'd829, 10'd830, 10'd831, 10'd832, 10'd833, 10'd834, 10'd835, 10'd836, 10'd837, 10'd838, 10'd839, 10'd840, 10'd841, 10'd842, 10'd843, 10'd844, 10'd845, 10'd846, 10'd847, 10'd848, 10'd849, 10'd850, 10'd851, 10'd852, 10'd853, 10'd854, 10'd855, 10'd856, 10'd857, 10'd858, 10'd859, 10'd860, 10'd861, 10'd862: sample = 3;
            10'd863, 10'd864, 10'd865, 10'd866, 10'd867, 10'd868, 10'd869, 10'd870, 10'd871, 10'd872, 10'd873, 10'd874, 10'd875, 10'd876, 10'd877, 10'd878, 10'd879, 10'd880, 10'd881, 10'd882, 10'd883, 10'd884, 10'd885, 10'd886, 10'd887, 10'd888, 10'd889, 10'd890, 10'd891, 10'd892, 10'd893, 10'd894, 10'd895, 10'd896, 10'd897, 10'd898, 10'd899, 10'd900, 10'd901, 10'd902, 10'd903, 10'd904, 10'd905, 10'd906, 10'd907, 10'd908, 10'd909, 10'd910, 10'd911, 10'd912, 10'd913, 10'd914, 10'd915, 10'd916, 10'd917, 10'd918, 10'd919: sample = 4;
            10'd920, 10'd921, 10'd922, 10'd923, 10'd924, 10'd925, 10'd926, 10'd927, 10'd928, 10'd929, 10'd930, 10'd931, 10'd932, 10'd933, 10'd934, 10'd935, 10'd936, 10'd937, 10'd938, 10'd939, 10'd940, 10'd941, 10'd942, 10'd943, 10'd944, 10'd945, 10'd946, 10'd947, 10'd948, 10'd949, 10'd950, 10'd951, 10'd952, 10'd953, 10'd954, 10'd955, 10'd956: sample = 5;
            10'd957, 10'd958, 10'd959, 10'd960, 10'd961, 10'd962, 10'd963, 10'd964, 10'd965, 10'd966, 10'd967, 10'd968, 10'd969, 10'd970, 10'd971, 10'd972, 10'd973, 10'd974, 10'd975, 10'd976, 10'd977: sample = 6;
            10'd978, 10'd979, 10'd980, 10'd981, 10'd982, 10'd983, 10'd984, 10'd985, 10'd986, 10'd987, 10'd988: sample = 7;
            10'd989, 10'd990, 10'd991, 10'd992, 10'd993: sample = 8;
            10'd994, 10'd995: sample = 9;
            10'd996: sample = 10;